module top_module(
    output zero
);// Module body starts after semicolon
    // Problem Statement 
    // Build a circuit with no inputs and one output that is constant LOW or ZERO
assign zero = 0;
    
endmodule
