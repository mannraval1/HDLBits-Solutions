module top_module( output one );
// Problem Statement
// Build a circuit with no inputs and outputs
// The output of the circuit should always drive 1 or HIGH logic
// Insert your code here
    assign one = 1'b1;

endmodule
